module inputs (
  input wire [0:7] data_i,
  input wire [0:7] mask_i,
  output wire [0:1] i_0,
  output wire [0:1] i_1,
  output wire [0:1] i_2,
  output wire [0:1] i_3,
  output wire [0:1] i_4,
  output wire [0:1] i_5, 
  output wire [0:1] i_6,
  output wire [0:1] i_7
);
  assign i_0[0:1] = { data_i[0], mask_i[0] };
  assign i_1[0:1] = { data_i[1], mask_i[1] };
  assign i_2[0:1] = { data_i[2], mask_i[2] };
  assign i_3[0:1] = { data_i[3], mask_i[3] };
  assign i_4[0:1] = { data_i[4], mask_i[4] };
  assign i_5[0:1] = { data_i[5], mask_i[5] };
  assign i_6[0:1] = { data_i[6], mask_i[6] };
  assign i_7[0:1] = { data_i[7], mask_i[7] };
endmodule


module outputs (
  input wire [0:7] data_o,
  input wire [0:7] mask_o,
  output wire [0:1] o_0,
  output wire [0:1] o_1,
  output wire [0:1] o_2,
  output wire [0:1] o_3,
  output wire [0:1] o_4,
  output wire [0:1] o_5,
  output wire [0:1] o_6,
  output wire [0:1] o_7
); 
  assign o_0[0:1] = { data_o[0], mask_o[0] };
  assign o_1[0:1] = { data_o[1], mask_o[1] };
  assign o_2[0:1] = { data_o[2], mask_o[2] };
  assign o_3[0:1] = { data_o[3], mask_o[3] };
  assign o_4[0:1] = { data_o[4], mask_o[4] };
  assign o_5[0:1] = { data_o[5], mask_o[5] };
  assign o_6[0:1] = { data_o[6], mask_o[6] };
  assign o_7[0:1] = { data_o[7], mask_o[7] };
endmodule


module randoms(
  input wire [0:27] prd_i,
  output wire [0:27] prd_in
);
  assign prd_in[0:27] = prd_i[0:27];
endmodule


module public_inputs(
  input wire clk_i,
  input wire rst_ni,
  input wire en_i,
  input wire out_ack_i,
  input [0:1] op_i,
  input [0:1] count_q_i,
  output wire clk_in,
  output wire rst_nin,
  output wire en_in,
  output wire out_ack_in,
  output wire op_i_0,
  output wire op_i_1,
  output wire count_q_i_0,
  output wire count_q_i_1
);
  assign clk_in = clk_i;
  assign rst_nin = rst_ni;
  assign en_in = en_i;
  assign out_ack_in = out_ack_i;
  assign op_i_0 = op_i[0];
  assign op_i_1 = op_i[1];
  assign count_q_i_0 = count_q_i[0];
  assign count_q_i_1 = count_q_i[1];
endmodule


module others(
  input wire out_req_o,
  input wire [0:19] prd_o,
  output wire out_req_out,
  output wire prd_o_0,
  output wire prd_o_1,
  output wire prd_o_2,
  output wire prd_o_3,
  output wire prd_o_4,
  output wire prd_o_5,
  output wire prd_o_6,
  output wire prd_o_7,
  output wire prd_o_8,
  output wire prd_o_9,
  output wire prd_o_10,
  output wire prd_o_11,
  output wire prd_o_12,
  output wire prd_o_13,
  output wire prd_o_14,
  output wire prd_o_15,
  output wire prd_o_16,
  output wire prd_o_17,
  output wire prd_o_18,
  output wire prd_o_19,
);
  assign out_req_out = out_req_o;
  assign prd_o_0 = prd_o[0];
  assign prd_o_1 = prd_o[1];
  assign prd_o_2 = prd_o[2];
  assign prd_o_3 = prd_o[3];
  assign prd_o_4 = prd_o[4];
  assign prd_o_5 = prd_o[5];
  assign prd_o_6 = prd_o[6];
  assign prd_o_7 = prd_o[7];
  assign prd_o_8 = prd_o[8];
  assign prd_o_9 = prd_o[9];
  assign prd_o_10 = prd_o[10];
  assign prd_o_11 = prd_o[11];
  assign prd_o_12 = prd_o[12];
  assign prd_o_13 = prd_o[13];
  assign prd_o_14 = prd_o[14];
  assign prd_o_15 = prd_o[15];
  assign prd_o_16 = prd_o[16];
  assign prd_o_17 = prd_o[17];
  assign prd_o_18 = prd_o[18];
  assign prd_o_19 = prd_o[19];

endmodule

