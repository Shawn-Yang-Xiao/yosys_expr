module aes_control_fsm_n (
	clk_i,
	rst_ni,
	ctrl_qe_i,
	ctrl_we_o,
	ctrl_phase_i,
	ctrl_err_storage_i,
	op_i,
	mode_i,
	cipher_op_i,
	sideload_i,
	prng_reseed_rate_i,
	manual_operation_i,
	key_touch_forces_reseed_i,
	start_i,
	key_iv_data_in_clear_i,
	data_out_clear_i,
	prng_reseed_i,
	mux_sel_err_i,
	sp_enc_err_i,
	lc_escalate_en_i,
	alert_fatal_i,
	alert_o,
	key_sideload_valid_i,
	key_init_qe_i,
	iv_qe_i,
	data_in_qe_i,
	data_out_re_i,
	data_in_we_o,
	data_out_we_no,
	data_in_prev_sel_o,
	data_in_prev_we_no,
	state_in_sel_o,
	add_state_in_sel_o,
	add_state_out_sel_o,
	ctr_incr_no,
	ctr_ready_ni,
	ctr_we_ni,
	cipher_in_valid_no,
	cipher_in_ready_ni,
	cipher_out_valid_ni,
	cipher_out_ready_no,
	cipher_crypt_no,
	cipher_crypt_ni,
	cipher_dec_key_gen_no,
	cipher_dec_key_gen_ni,
	cipher_prng_reseed_o,
	cipher_prng_reseed_i,
	cipher_key_clear_o,
	cipher_key_clear_i,
	cipher_data_out_clear_o,
	cipher_data_out_clear_i,
	key_init_sel_o,
	key_init_we_no,
	iv_sel_o,
	iv_we_no,
	prng_data_req_o,
	prng_data_ack_i,
	prng_reseed_req_o,
	prng_reseed_ack_i,
	start_we_o,
	key_iv_data_in_clear_we_o,
	data_out_clear_we_o,
	prng_reseed_o,
	prng_reseed_we_o,
	idle_o,
	idle_we_o,
	stall_o,
	stall_we_o,
	output_lost_i,
	output_lost_o,
	output_lost_we_o,
	output_valid_o,
	output_valid_we_o,
	input_ready_o,
	input_ready_we_o
);
	parameter [0:0] SecMasking = 0;
	input wire clk_i;
	input wire rst_ni;
	input wire ctrl_qe_i;
	output wire ctrl_we_o;
	input wire ctrl_phase_i;
	input wire ctrl_err_storage_i;
	localparam signed [31:0] aes_pkg_AES_OP_WIDTH = 2;
	input wire [1:0] op_i;
	localparam signed [31:0] aes_pkg_AES_MODE_WIDTH = 6;
	input wire [5:0] mode_i;
	input wire [1:0] cipher_op_i;
	input wire sideload_i;
	localparam signed [31:0] aes_pkg_AES_PRNGRESEEDRATE_WIDTH = 3;
	input wire [2:0] prng_reseed_rate_i;
	input wire manual_operation_i;
	input wire key_touch_forces_reseed_i;
	input wire start_i;
	input wire key_iv_data_in_clear_i;
	input wire data_out_clear_i;
	input wire prng_reseed_i;
	input wire mux_sel_err_i;
	input wire sp_enc_err_i;
	localparam signed [31:0] lc_ctrl_pkg_TxWidth = 4;
	input wire [3:0] lc_escalate_en_i;
	input wire alert_fatal_i;
	output wire alert_o;
	input wire key_sideload_valid_i;
	localparam [31:0] aes_pkg_NumSharesKey = 2;
	localparam signed [31:0] aes_reg_pkg_NumRegsKey = 8;
	input wire [(aes_pkg_NumSharesKey * aes_reg_pkg_NumRegsKey) - 1:0] key_init_qe_i;
	localparam signed [31:0] aes_reg_pkg_NumRegsIv = 4;
	input wire [3:0] iv_qe_i;
	localparam signed [31:0] aes_reg_pkg_NumRegsData = 4;
	input wire [3:0] data_in_qe_i;
	input wire [3:0] data_out_re_i;
	output wire data_in_we_o;
	output wire data_out_we_no;
	localparam signed [31:0] aes_pkg_Mux2SelWidth = 3;
	localparam signed [31:0] aes_pkg_DIPSelWidth = aes_pkg_Mux2SelWidth;
	output wire [2:0] data_in_prev_sel_o;
	output wire data_in_prev_we_no;
	localparam signed [31:0] aes_pkg_SISelWidth = aes_pkg_Mux2SelWidth;
	output wire [2:0] state_in_sel_o;
	localparam signed [31:0] aes_pkg_AddSISelWidth = aes_pkg_Mux2SelWidth;
	output wire [2:0] add_state_in_sel_o;
	localparam signed [31:0] aes_pkg_Mux3SelWidth = 5;
	localparam signed [31:0] aes_pkg_AddSOSelWidth = aes_pkg_Mux3SelWidth;
	output wire [4:0] add_state_out_sel_o;
	output wire ctr_incr_no;
	input wire ctr_ready_ni;
	localparam [31:0] aes_pkg_SliceSizeCtr = 16;
	localparam [31:0] aes_pkg_NumSlicesCtr = 8;
	input wire [7:0] ctr_we_ni;
	output wire cipher_in_valid_no;
	input wire cipher_in_ready_ni;
	input wire cipher_out_valid_ni;
	output wire cipher_out_ready_no;
	output wire cipher_crypt_no;
	input wire cipher_crypt_ni;
	output wire cipher_dec_key_gen_no;
	input wire cipher_dec_key_gen_ni;
	output wire cipher_prng_reseed_o;
	input wire cipher_prng_reseed_i;
	output wire cipher_key_clear_o;
	input wire cipher_key_clear_i;
	output wire cipher_data_out_clear_o;
	input wire cipher_data_out_clear_i;
	localparam signed [31:0] aes_pkg_KeyInitSelWidth = aes_pkg_Mux3SelWidth;
	output wire [4:0] key_init_sel_o;
	output wire [(aes_pkg_NumSharesKey * aes_reg_pkg_NumRegsKey) - 1:0] key_init_we_no;
	localparam signed [31:0] aes_pkg_Mux6SelWidth = 6;
	localparam signed [31:0] aes_pkg_IVSelWidth = aes_pkg_Mux6SelWidth;
	output wire [5:0] iv_sel_o;
	output wire [7:0] iv_we_no;
	output wire prng_data_req_o;
	input wire prng_data_ack_i;
	output wire prng_reseed_req_o;
	input wire prng_reseed_ack_i;
	output wire start_we_o;
	output wire key_iv_data_in_clear_we_o;
	output wire data_out_clear_we_o;
	output wire prng_reseed_o;
	output wire prng_reseed_we_o;
	output wire idle_o;
	output wire idle_we_o;
	output wire stall_o;
	output wire stall_we_o;
	input wire output_lost_i;
	output wire output_lost_o;
	output wire output_lost_we_o;
	output wire output_valid_o;
	output wire output_valid_we_o;
	output wire input_ready_o;
	output wire input_ready_we_o;
	localparam signed [31:0] NumInBufBits = ((((((31 + (aes_pkg_NumSharesKey * aes_reg_pkg_NumRegsKey)) + aes_reg_pkg_NumRegsIv) + aes_reg_pkg_NumRegsData) + aes_reg_pkg_NumRegsData) + 1) + aes_pkg_NumSlicesCtr) + 10;
	wire [NumInBufBits - 1:0] in;
	wire [NumInBufBits - 1:0] in_buf;
	assign in = {ctrl_qe_i, ctrl_phase_i, ctrl_err_storage_i, op_i, mode_i, cipher_op_i, sideload_i, prng_reseed_rate_i, manual_operation_i, key_touch_forces_reseed_i, start_i, key_iv_data_in_clear_i, data_out_clear_i, prng_reseed_i, mux_sel_err_i, sp_enc_err_i, lc_escalate_en_i, alert_fatal_i, key_sideload_valid_i, key_init_qe_i, iv_qe_i, data_in_qe_i, data_out_re_i, ctr_ready_ni, ctr_we_ni, cipher_in_ready_ni, cipher_out_valid_ni, cipher_crypt_ni, cipher_dec_key_gen_ni, cipher_prng_reseed_i, cipher_key_clear_i, cipher_data_out_clear_i, prng_data_ack_i, prng_reseed_ack_i, output_lost_i};
	prim_xilinx_buf #(.Width(NumInBufBits)) u_prim_xilinx_buf_in(
		.in_i(in),
		.out_o(in_buf)
	);
	wire ctrl_qe;
	wire ctrl_phase;
	wire ctrl_err_storage;
	wire [1:0] op;
	wire [5:0] mode;
	wire [1:0] cipher_op;
	wire [1:0] cipher_op_raw;
	wire sideload;
	wire [2:0] prng_reseed_rate;
	wire manual_operation;
	wire key_touch_forces_reseed;
	wire start;
	wire key_iv_data_in_clear;
	wire data_out_clear;
	wire prng_reseed_in_buf;
	wire mux_sel_err;
	wire sp_enc_err;
	wire [3:0] lc_escalate_en;
	wire alert_fatal;
	wire key_sideload_valid;
	wire [(aes_pkg_NumSharesKey * aes_reg_pkg_NumRegsKey) - 1:0] key_init_qe;
	wire [3:0] iv_qe;
	wire [3:0] data_in_qe;
	wire [3:0] data_out_re;
	wire ctr_ready_n;
	wire [7:0] ctr_we_n;
	wire cipher_in_ready_n;
	wire cipher_out_valid_n;
	wire cipher_crypt_in_buf_n;
	wire cipher_dec_key_gen_in_buf_n;
	wire cipher_prng_reseed_in_buf;
	wire cipher_key_clear_in_buf;
	wire cipher_data_out_clear_in_buf;
	wire prng_data_ack;
	wire prng_reseed_ack;
	wire output_lost_in_buf;
	assign {ctrl_qe, ctrl_phase, ctrl_err_storage, op, mode, cipher_op_raw, sideload, prng_reseed_rate, manual_operation, key_touch_forces_reseed, start, key_iv_data_in_clear, data_out_clear, prng_reseed_in_buf, mux_sel_err, sp_enc_err, lc_escalate_en, alert_fatal, key_sideload_valid, key_init_qe, iv_qe, data_in_qe, data_out_re, ctr_ready_n, ctr_we_n, cipher_in_ready_n, cipher_out_valid_n, cipher_crypt_in_buf_n, cipher_dec_key_gen_in_buf_n, cipher_prng_reseed_in_buf, cipher_key_clear_in_buf, cipher_data_out_clear_in_buf, prng_data_ack, prng_reseed_ack, output_lost_in_buf} = in_buf;
	function automatic [1:0] sv2v_cast_E41EB;
		input reg [1:0] inp;
		sv2v_cast_E41EB = inp;
	endfunction
	assign cipher_op = sv2v_cast_E41EB(cipher_op_raw);
	wire ctrl_we;
	wire alert;
	wire data_in_we;
	wire data_out_we;
	wire [2:0] data_in_prev_sel;
	wire data_in_prev_we;
	wire [2:0] state_in_sel;
	wire [2:0] add_state_in_sel;
	wire [4:0] add_state_out_sel;
	wire ctr_incr;
	wire cipher_in_valid;
	wire cipher_out_ready;
	wire cipher_crypt_out_buf;
	wire cipher_dec_key_gen_out_buf;
	wire cipher_prng_reseed_out_buf;
	wire cipher_key_clear_out_buf;
	wire cipher_data_out_clear_out_buf;
	wire [4:0] key_init_sel;
	wire [(aes_pkg_NumSharesKey * aes_reg_pkg_NumRegsKey) - 1:0] key_init_we;
	wire [5:0] iv_sel;
	wire [7:0] iv_we;
	wire prng_data_req;
	wire prng_reseed_req;
	wire start_we;
	wire key_iv_data_in_clear_we;
	wire data_out_clear_we;
	wire prng_reseed_out_buf;
	wire prng_reseed_we;
	wire idle;
	wire idle_we;
	wire stall;
	wire stall_we;
	wire output_lost_out_buf;
	wire output_lost_we;
	wire output_valid;
	wire output_valid_we;
	wire input_ready;
	wire input_ready_we;
	aes_control_fsm #(.SecMasking(SecMasking)) u_aes_control_fsm(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.ctrl_qe_i(ctrl_qe),
		.ctrl_we_o(ctrl_we),
		.ctrl_phase_i(ctrl_phase),
		.ctrl_err_storage_i(ctrl_err_storage),
		.op_i(op),
		.mode_i(mode),
		.cipher_op_i(cipher_op),
		.sideload_i(sideload),
		.prng_reseed_rate_i(prng_reseed_rate),
		.manual_operation_i(manual_operation),
		.key_touch_forces_reseed_i(key_touch_forces_reseed),
		.start_i(start),
		.key_iv_data_in_clear_i(key_iv_data_in_clear),
		.data_out_clear_i(data_out_clear),
		.prng_reseed_i(prng_reseed_in_buf),
		.mux_sel_err_i(mux_sel_err),
		.sp_enc_err_i(sp_enc_err),
		.lc_escalate_en_i(lc_escalate_en),
		.alert_fatal_i(alert_fatal),
		.alert_o(alert),
		.key_sideload_valid_i(key_sideload_valid),
		.key_init_qe_i(key_init_qe),
		.iv_qe_i(iv_qe),
		.data_in_qe_i(data_in_qe),
		.data_out_re_i(data_out_re),
		.data_in_we_o(data_in_we),
		.data_out_we_o(data_out_we),
		.data_in_prev_sel_o(data_in_prev_sel),
		.data_in_prev_we_o(data_in_prev_we),
		.state_in_sel_o(state_in_sel),
		.add_state_in_sel_o(add_state_in_sel),
		.add_state_out_sel_o(add_state_out_sel),
		.ctr_incr_o(ctr_incr),
		.ctr_ready_i(~ctr_ready_n),
		.ctr_we_i(~ctr_we_n),
		.cipher_in_valid_o(cipher_in_valid),
		.cipher_in_ready_i(~cipher_in_ready_n),
		.cipher_out_valid_i(~cipher_out_valid_n),
		.cipher_out_ready_o(cipher_out_ready),
		.cipher_crypt_o(cipher_crypt_out_buf),
		.cipher_crypt_i(~cipher_crypt_in_buf_n),
		.cipher_dec_key_gen_o(cipher_dec_key_gen_out_buf),
		.cipher_dec_key_gen_i(~cipher_dec_key_gen_in_buf_n),
		.cipher_prng_reseed_o(cipher_prng_reseed_out_buf),
		.cipher_prng_reseed_i(cipher_prng_reseed_in_buf),
		.cipher_key_clear_o(cipher_key_clear_out_buf),
		.cipher_key_clear_i(cipher_key_clear_in_buf),
		.cipher_data_out_clear_o(cipher_data_out_clear_out_buf),
		.cipher_data_out_clear_i(cipher_data_out_clear_in_buf),
		.key_init_sel_o(key_init_sel),
		.key_init_we_o(key_init_we),
		.iv_sel_o(iv_sel),
		.iv_we_o(iv_we),
		.prng_data_req_o(prng_data_req),
		.prng_data_ack_i(prng_data_ack),
		.prng_reseed_req_o(prng_reseed_req),
		.prng_reseed_ack_i(prng_reseed_ack),
		.start_we_o(start_we),
		.key_iv_data_in_clear_we_o(key_iv_data_in_clear_we),
		.data_out_clear_we_o(data_out_clear_we),
		.prng_reseed_o(prng_reseed_out_buf),
		.prng_reseed_we_o(prng_reseed_we),
		.idle_o(idle),
		.idle_we_o(idle_we),
		.stall_o(stall),
		.stall_we_o(stall_we),
		.output_lost_i(output_lost_in_buf),
		.output_lost_o(output_lost_out_buf),
		.output_lost_we_o(output_lost_we),
		.output_valid_o(output_valid),
		.output_valid_we_o(output_valid_we),
		.input_ready_o(input_ready),
		.input_ready_we_o(input_ready_we)
	);
	localparam signed [31:0] NumOutBufBits = (((32 + (aes_pkg_NumSharesKey * aes_reg_pkg_NumRegsKey)) + aes_pkg_IVSelWidth) + aes_pkg_NumSlicesCtr) + 17;
	wire [NumOutBufBits - 1:0] out;
	wire [NumOutBufBits - 1:0] out_buf;
	assign out = {ctrl_we, alert, data_in_we, ~data_out_we, data_in_prev_sel, ~data_in_prev_we, state_in_sel, add_state_in_sel, add_state_out_sel, ~ctr_incr, ~cipher_in_valid, ~cipher_out_ready, ~cipher_crypt_out_buf, ~cipher_dec_key_gen_out_buf, cipher_prng_reseed_out_buf, cipher_key_clear_out_buf, cipher_data_out_clear_out_buf, key_init_sel, ~key_init_we, iv_sel, ~iv_we, prng_data_req, prng_reseed_req, start_we, key_iv_data_in_clear_we, data_out_clear_we, prng_reseed_out_buf, prng_reseed_we, idle, idle_we, stall, stall_we, output_lost_out_buf, output_lost_we, output_valid, output_valid_we, input_ready, input_ready_we};
	prim_xilinx_buf #(.Width(NumOutBufBits)) u_prim_xilinx_buf_out(
		.in_i(out),
		.out_o(out_buf)
	);
	assign {ctrl_we_o, alert_o, data_in_we_o, data_out_we_no, data_in_prev_sel_o, data_in_prev_we_no, state_in_sel_o, add_state_in_sel_o, add_state_out_sel_o, ctr_incr_no, cipher_in_valid_no, cipher_out_ready_no, cipher_crypt_no, cipher_dec_key_gen_no, cipher_prng_reseed_o, cipher_key_clear_o, cipher_data_out_clear_o, key_init_sel_o, key_init_we_no, iv_sel_o, iv_we_no, prng_data_req_o, prng_reseed_req_o, start_we_o, key_iv_data_in_clear_we_o, data_out_clear_we_o, prng_reseed_o, prng_reseed_we_o, idle_o, idle_we_o, stall_o, stall_we_o, output_lost_o, output_lost_we_o, output_valid_o, output_valid_we_o, input_ready_o, input_ready_we_o} = out_buf;
endmodule
